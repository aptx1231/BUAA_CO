`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:53:56 11/24/2018 
// Design Name: 
// Module Name:    controller 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module controller(
	 input [5:0] op,
	 input [5:0] func,
	 input [4:0] rt,
    output reg[3:0] ALUCtrl,
    output reg[1:0] RegDst,
    output reg ALUASrc,
	 output reg ALUBSrc,
    output reg RegWrite,
    output reg MemRead,
    output reg MemWrite,
    output reg [1:0] MemtoReg,
    output reg [1:0]ExtOp,
    output reg if_beq,
	 output reg if_bne,
	 output reg if_blez,
	 output reg if_bgez,
	 output reg if_bltz,
	 output reg if_bgtz,
    output reg if_j,
	 output reg [1:0]PCsel,
	 output reg if_sh,
	 output reg if_sb,
	 output reg[2:0] dataOp,
	 output reg[1:0] multdivOp,
	 output reg start,
	 output reg if_mthi,
	 output reg if_mtlo,
	 output reg if_mfhi,
	 output reg if_mflo
    );
	 initial  begin
		PCsel <= 2'b00;
	 end
	always@(*) 
	begin
		case (op)
		6'b000000://R 
		begin
			RegDst<=2'b01;
			ALUBSrc<=0;
			MemRead<=0;
			MemWrite<=0;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			if_sh<=0;
			if_sb<=0;
			if_j<=0;
			dataOp<=3'b000;
			case(func)
				6'b100001: begin  //addu
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0010;
					PCsel<=2'b00;	
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b100000: begin  //add
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0010;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b100011: begin  //subu
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0011;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b100010: begin  //sub
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0011;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b100100: begin  //and
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0000;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b100101: begin  //or
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0001;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b100110: begin  //xor
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0100;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b100111: begin  //nor
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0101;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b001000: begin  //jr
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0000;
					PCsel<=2'b01;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b001001: begin  //jalr
					ALUASrc<=0;
					MemtoReg<=2'b10;
					ALUCtrl<=4'b0000;
					PCsel<=2'b01;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b000000: begin  //sll nop
					ALUASrc<=1;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0110;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b000100: begin  //sllv
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0110;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b000010: begin  //srl
					ALUASrc<=1;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0111;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b000110: begin  //srlv
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0111;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b000011: begin  //sra
					ALUASrc<=1;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b1000;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b000111: begin  //srav
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b1000;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b101010: begin  //slt
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b1001;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b101011: begin  //sltu
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b1010;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b011000: begin  //mult
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0000;
					PCsel<=2'b00;
					RegWrite<=0;
					multdivOp<=2'b00;		
					start<=1;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b011001: begin  //multu
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0000;
					PCsel<=2'b00;
					RegWrite<=0;	
					multdivOp<=2'b01;
					start<=1;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b011010: begin  //div
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0000;
					PCsel<=2'b00;
					RegWrite<=0;
					multdivOp<=2'b10;		
					start<=1;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b011011: begin  //divu
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0000;
					PCsel<=2'b00;
					RegWrite<=0;	
					multdivOp<=2'b11;
					start<=1;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b010000: begin  //mfhi
					ALUASrc<=0;
					MemtoReg<=2'b11;
					ALUCtrl<=4'b0000;
					PCsel<=2'b00;
					RegWrite<=1;
					multdivOp<=2'b00;		
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=1;
					if_mflo<=0;
				end
				6'b010010: begin  //mflo
					ALUASrc<=0;
					MemtoReg<=2'b11;
					ALUCtrl<=4'b0000;
					PCsel<=2'b00;
					RegWrite<=1;	
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=1;
				end
				6'b010001: begin  //mthi
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0000;
					PCsel<=2'b00;
					RegWrite<=0;
					multdivOp<=2'b00;		
					start<=0;
					if_mthi<=1;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
				end
				6'b010011: begin  //mtlo
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0000;
					PCsel<=2'b00;
					RegWrite<=0;	
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=1;
					if_mfhi<=0;
					if_mflo<=0;
				end
				default:  begin
					ALUASrc<=0;
					MemtoReg<=2'b00;
					ALUCtrl<=4'b0000;
					PCsel<=2'b00;
					RegWrite<=1;	
					multdivOp<=2'b00;
					start<=0;
					if_mthi<=0;
					if_mtlo<=0;
					if_mfhi<=0;
					if_mflo<=0;
					end
			endcase
		end
		6'b100011://lw
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=1;
			MemWrite<=0;
			MemtoReg<=2'b01;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b100000://lb
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=1;
			MemWrite<=0;
			MemtoReg<=2'b01;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b010;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b100100://lbu
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=1;
			MemWrite<=0;
			MemtoReg<=2'b01;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b001;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b100001://lh
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=1;
			MemWrite<=0;
			MemtoReg<=2'b01;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b100;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b100101://lhb
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=1;
			MemWrite<=0;
			MemtoReg<=2'b01;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b011;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b101011://sw
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=0;
			MemRead<=0;
			MemWrite<=1;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b101001://sh
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=0;
			MemRead<=0;
			MemWrite<=1;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=1;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b101000://sb
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=0;
			MemRead<=0;
			MemWrite<=1;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=1;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
      6'b000100://beq
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=0;
			RegWrite<=0;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=1;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0000;
			if_j<=0;
			PCsel<=2'b10;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;	
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;		
		end
		
		6'b000101://bne
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=0;
			RegWrite<=0;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=1;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0000;
			if_j<=0;
			PCsel<=2'b10;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
 
		6'b000111://bgtz
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=0;
			RegWrite<=0;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=1;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0000;
			if_j<=0;
			PCsel<=2'b10;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b000110://blez
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=0;
			RegWrite<=0;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=1;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0000;
			if_j<=0;
			PCsel<=2'b10;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b000001://bgez/bltz
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=0;
			RegWrite<=0;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			ALUCtrl<=4'b0000;
			if_j<=0;
			PCsel<=2'b10;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
			case(rt) 
				5'b00001:begin//bgez
					if_bgez<=1;
					if_bltz<=0;
				end
				5'b00000:begin//bltz
					if_bgez<=0;
					if_bltz<=1;
				end
				default:begin
					if_bgez<=0;
					if_bltz<=0;
				end
			endcase
		end
		
      6'b001111://lui
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b10;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end

      6'b001101://ori
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b01;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0001;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b001010://slti
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b1001;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b001011://sltiu
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b1010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b001100://andi
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b01;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0000;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b001110://xori
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b01;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0100;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b001001://addiu
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end

		6'b001000://addi
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=1;
			RegWrite<=1;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0010;
			if_j<=0;
			PCsel<=2'b00;
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b000011://jal
		begin
			RegDst<=2'b10;
			ALUASrc<=0;
			ALUBSrc<=0;
			RegWrite<=1;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b10;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0000;
			if_j<=1;
			PCsel<=2'b10;	
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		
		6'b000010://j
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=0;
			RegWrite<=0;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0000;
			if_j<=1;
			PCsel<=2'b10;	
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end

		default: 
		begin
			RegDst<=2'b00;
			ALUASrc<=0;
			ALUBSrc<=0;
			RegWrite<=0;
			MemRead<=0;
			MemWrite<=0;
			MemtoReg<=2'b00;
			ExtOp<=2'b00;
			if_beq<=0;
			if_bne<=0;
			if_bgtz<=0;
			if_blez<=0;
			if_bgez<=0;
			if_bltz<=0;
			ALUCtrl<=4'b0000;
			if_j<=0;
			PCsel<=2'b00;	
			if_sh<=0;
			if_sb<=0;
			dataOp<=3'b000;
			multdivOp<=2'b00;
			start<=0;
			if_mthi<=0;
			if_mtlo<=0;
			if_mfhi<=0;
			if_mflo<=0;
		end
		endcase
	end	

endmodule
